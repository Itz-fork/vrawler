module huvl