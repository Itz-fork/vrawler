module vrawler