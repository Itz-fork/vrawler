module huv